interface SPI_IF(clk);
 logic MOSI,rst_n,SS_n,MISO;
 logic [2:0] dut_state;
 input clk;
	
endinterface : SPI_IF